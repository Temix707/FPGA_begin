library verilog;
use verilog.vl_types.all;
entity lab5_vlg_vec_tst is
end lab5_vlg_vec_tst;
