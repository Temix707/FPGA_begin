library verilog;
use verilog.vl_types.all;
entity lr4dop_vlg_vec_tst is
end lr4dop_vlg_vec_tst;
