library verilog;
use verilog.vl_types.all;
entity check_me_1_vlg_vec_tst is
end check_me_1_vlg_vec_tst;
