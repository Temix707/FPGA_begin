library verilog;
use verilog.vl_types.all;
entity lr6_vlg_vec_tst is
end lr6_vlg_vec_tst;
