/*module shift_reg_out_l4(

	input CLOCK_50,
	input [1:0] KEY,
	input [0:0]SW,
	//input ISL, 
	
	//output OSL,
	output [9:0] LEDR,
	output [6:0] HEX0

);


shift_reg_l4 init_1 (CLOCK_50, KEY[1:0], SW[0:0], LEDR[9:0], HEX0[6:0]);



endmodule
*/